//dummy wrapper of xilinx fifo, replace your code here

module wstrb_fifo (
);

endmodule
