//dummy wrapper of xilinx fifo, replace your code here

module rdata_fifo (
);


endmodule
