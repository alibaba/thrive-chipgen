//dummy wrapper of xilinx fifo, replace your code here

module rinfo_fifo (
);

endmodule
