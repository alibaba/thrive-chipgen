//dummy wrapper of xilinx fifo, replace your code here

module wdata_fifo (
);

endmodule
