//dummy wrapper of xilinx fifo, replace your code here

module wcmd_fifo (
);

endmodule