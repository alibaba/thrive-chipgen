/* 
*Copyright (c) 2021, Alibaba Group;
*Licensed under the Apache License, Version 2.0 (the "License");
*you may not use this file except in compliance with the License.
*You may obtain a copy of the License at

*   http://www.apache.org/licenses/LICENSE-2.0

*Unless required by applicable law or agreed to in writing, software
*distributed under the License is distributed on an "AS IS" BASIS,
*WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
*See the License for the specific language governing permissions and
*limitations under the License.
*/

// Dumping Control
`ifndef NO_DUMP
initial
begin
    `ifdef VCS
        $fsdbAutoSwitchDumpfile(3000,"top_debug.fsdb",3);
        $fsdbDumpvars(0, tb_top, "+mda");
    `else
        $dumpfile("top_debug.vcd");
        $dumpvars();
    `endif//VCS
end
`endif//NO_DUMP
